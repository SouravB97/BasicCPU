`define ADDB 'h00 //ADD B to Ac and store in Ac
