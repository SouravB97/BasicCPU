`define ADDB 'h02 //ADD B to Ac and store in Ac
