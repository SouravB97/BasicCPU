`define ADDB 'h02 //ADD B to Ac and store in Ac
`define ANDB 'h08 //AND B to Ac and store in Ac
